/*
    
*/
module test;
endmodule 